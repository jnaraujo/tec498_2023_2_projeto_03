module projeto();

endmodule
